// system_acl_iface_acl_kernel_interface.v

// Generated using ACDS version 14.1 186 at 2023.12.14.11:25:57

`timescale 1 ps / 1 ps
module system_acl_iface_acl_kernel_interface (
		input  wire        clk_clk,                    //                    clk.clk
		input  wire        reset_reset_n,              //                  reset.reset_n
		output wire        kernel_cntrl_waitrequest,   //           kernel_cntrl.waitrequest
		output wire [31:0] kernel_cntrl_readdata,      //                       .readdata
		output wire        kernel_cntrl_readdatavalid, //                       .readdatavalid
		input  wire [0:0]  kernel_cntrl_burstcount,    //                       .burstcount
		input  wire [31:0] kernel_cntrl_writedata,     //                       .writedata
		input  wire [13:0] kernel_cntrl_address,       //                       .address
		input  wire        kernel_cntrl_write,         //                       .write
		input  wire        kernel_cntrl_read,          //                       .read
		input  wire [3:0]  kernel_cntrl_byteenable,    //                       .byteenable
		input  wire        kernel_cntrl_debugaccess,   //                       .debugaccess
		input  wire        kernel_cra_waitrequest,     //             kernel_cra.waitrequest
		input  wire [63:0] kernel_cra_readdata,        //                       .readdata
		input  wire        kernel_cra_readdatavalid,   //                       .readdatavalid
		output wire [0:0]  kernel_cra_burstcount,      //                       .burstcount
		output wire [63:0] kernel_cra_writedata,       //                       .writedata
		output wire [29:0] kernel_cra_address,         //                       .address
		output wire        kernel_cra_write,           //                       .write
		output wire        kernel_cra_read,            //                       .read
		output wire [7:0]  kernel_cra_byteenable,      //                       .byteenable
		output wire        kernel_cra_debugaccess,     //                       .debugaccess
		input  wire [0:0]  kernel_irq_from_kernel_irq, // kernel_irq_from_kernel.irq
		output wire [1:0]  acl_bsp_memorg_kernel_mode, //  acl_bsp_memorg_kernel.mode
		output wire [1:0]  acl_bsp_memorg_host_mode,   //    acl_bsp_memorg_host.mode
		input  wire        sw_reset_in_reset,          //            sw_reset_in.reset
		input  wire        kernel_clk_clk,             //             kernel_clk.clk
		output wire        sw_reset_export_reset_n,    //        sw_reset_export.reset_n
		output wire        kernel_reset_reset_n,       //           kernel_reset.reset_n
		output wire        kernel_irq_to_host_irq      //     kernel_irq_to_host.irq
	);

	wire         reset_controller_sw_reset_out_reset;                                    // reset_controller_sw:reset_out -> [irq_bridge_0:reset, kernel_cra:reset, mm_interconnect_0:kernel_cra_reset_reset_bridge_in_reset_reset, reset_controller_sw_reset_out_reset:in]
	wire         address_span_extender_0_expanded_master_waitrequest;                    // mm_interconnect_0:address_span_extender_0_expanded_master_waitrequest -> address_span_extender_0:avm_m0_waitrequest
	wire  [31:0] address_span_extender_0_expanded_master_readdata;                       // mm_interconnect_0:address_span_extender_0_expanded_master_readdata -> address_span_extender_0:avm_m0_readdata
	wire  [29:0] address_span_extender_0_expanded_master_address;                        // address_span_extender_0:avm_m0_address -> mm_interconnect_0:address_span_extender_0_expanded_master_address
	wire         address_span_extender_0_expanded_master_read;                           // address_span_extender_0:avm_m0_read -> mm_interconnect_0:address_span_extender_0_expanded_master_read
	wire   [3:0] address_span_extender_0_expanded_master_byteenable;                     // address_span_extender_0:avm_m0_byteenable -> mm_interconnect_0:address_span_extender_0_expanded_master_byteenable
	wire         address_span_extender_0_expanded_master_readdatavalid;                  // mm_interconnect_0:address_span_extender_0_expanded_master_readdatavalid -> address_span_extender_0:avm_m0_readdatavalid
	wire         address_span_extender_0_expanded_master_write;                          // address_span_extender_0:avm_m0_write -> mm_interconnect_0:address_span_extender_0_expanded_master_write
	wire  [31:0] address_span_extender_0_expanded_master_writedata;                      // address_span_extender_0:avm_m0_writedata -> mm_interconnect_0:address_span_extender_0_expanded_master_writedata
	wire   [0:0] address_span_extender_0_expanded_master_burstcount;                     // address_span_extender_0:avm_m0_burstcount -> mm_interconnect_0:address_span_extender_0_expanded_master_burstcount
	wire  [63:0] mm_interconnect_0_kernel_cra_s0_readdata;                               // kernel_cra:s0_readdata -> mm_interconnect_0:kernel_cra_s0_readdata
	wire         mm_interconnect_0_kernel_cra_s0_waitrequest;                            // kernel_cra:s0_waitrequest -> mm_interconnect_0:kernel_cra_s0_waitrequest
	wire         mm_interconnect_0_kernel_cra_s0_debugaccess;                            // mm_interconnect_0:kernel_cra_s0_debugaccess -> kernel_cra:s0_debugaccess
	wire  [29:0] mm_interconnect_0_kernel_cra_s0_address;                                // mm_interconnect_0:kernel_cra_s0_address -> kernel_cra:s0_address
	wire         mm_interconnect_0_kernel_cra_s0_read;                                   // mm_interconnect_0:kernel_cra_s0_read -> kernel_cra:s0_read
	wire   [7:0] mm_interconnect_0_kernel_cra_s0_byteenable;                             // mm_interconnect_0:kernel_cra_s0_byteenable -> kernel_cra:s0_byteenable
	wire         mm_interconnect_0_kernel_cra_s0_readdatavalid;                          // kernel_cra:s0_readdatavalid -> mm_interconnect_0:kernel_cra_s0_readdatavalid
	wire         mm_interconnect_0_kernel_cra_s0_write;                                  // mm_interconnect_0:kernel_cra_s0_write -> kernel_cra:s0_write
	wire  [63:0] mm_interconnect_0_kernel_cra_s0_writedata;                              // mm_interconnect_0:kernel_cra_s0_writedata -> kernel_cra:s0_writedata
	wire   [0:0] mm_interconnect_0_kernel_cra_s0_burstcount;                             // mm_interconnect_0:kernel_cra_s0_burstcount -> kernel_cra:s0_burstcount
	wire         kernel_cntrl_m0_waitrequest;                                            // mm_interconnect_1:kernel_cntrl_m0_waitrequest -> kernel_cntrl:m0_waitrequest
	wire  [31:0] kernel_cntrl_m0_readdata;                                               // mm_interconnect_1:kernel_cntrl_m0_readdata -> kernel_cntrl:m0_readdata
	wire         kernel_cntrl_m0_debugaccess;                                            // kernel_cntrl:m0_debugaccess -> mm_interconnect_1:kernel_cntrl_m0_debugaccess
	wire  [13:0] kernel_cntrl_m0_address;                                                // kernel_cntrl:m0_address -> mm_interconnect_1:kernel_cntrl_m0_address
	wire         kernel_cntrl_m0_read;                                                   // kernel_cntrl:m0_read -> mm_interconnect_1:kernel_cntrl_m0_read
	wire   [3:0] kernel_cntrl_m0_byteenable;                                             // kernel_cntrl:m0_byteenable -> mm_interconnect_1:kernel_cntrl_m0_byteenable
	wire         kernel_cntrl_m0_readdatavalid;                                          // mm_interconnect_1:kernel_cntrl_m0_readdatavalid -> kernel_cntrl:m0_readdatavalid
	wire  [31:0] kernel_cntrl_m0_writedata;                                              // kernel_cntrl:m0_writedata -> mm_interconnect_1:kernel_cntrl_m0_writedata
	wire         kernel_cntrl_m0_write;                                                  // kernel_cntrl:m0_write -> mm_interconnect_1:kernel_cntrl_m0_write
	wire   [0:0] kernel_cntrl_m0_burstcount;                                             // kernel_cntrl:m0_burstcount -> mm_interconnect_1:kernel_cntrl_m0_burstcount
	wire  [31:0] mm_interconnect_1_address_span_extender_0_windowed_slave_readdata;      // address_span_extender_0:avs_s0_readdata -> mm_interconnect_1:address_span_extender_0_windowed_slave_readdata
	wire         mm_interconnect_1_address_span_extender_0_windowed_slave_waitrequest;   // address_span_extender_0:avs_s0_waitrequest -> mm_interconnect_1:address_span_extender_0_windowed_slave_waitrequest
	wire   [9:0] mm_interconnect_1_address_span_extender_0_windowed_slave_address;       // mm_interconnect_1:address_span_extender_0_windowed_slave_address -> address_span_extender_0:avs_s0_address
	wire         mm_interconnect_1_address_span_extender_0_windowed_slave_read;          // mm_interconnect_1:address_span_extender_0_windowed_slave_read -> address_span_extender_0:avs_s0_read
	wire   [3:0] mm_interconnect_1_address_span_extender_0_windowed_slave_byteenable;    // mm_interconnect_1:address_span_extender_0_windowed_slave_byteenable -> address_span_extender_0:avs_s0_byteenable
	wire         mm_interconnect_1_address_span_extender_0_windowed_slave_readdatavalid; // address_span_extender_0:avs_s0_readdatavalid -> mm_interconnect_1:address_span_extender_0_windowed_slave_readdatavalid
	wire         mm_interconnect_1_address_span_extender_0_windowed_slave_write;         // mm_interconnect_1:address_span_extender_0_windowed_slave_write -> address_span_extender_0:avs_s0_write
	wire  [31:0] mm_interconnect_1_address_span_extender_0_windowed_slave_writedata;     // mm_interconnect_1:address_span_extender_0_windowed_slave_writedata -> address_span_extender_0:avs_s0_writedata
	wire   [0:0] mm_interconnect_1_address_span_extender_0_windowed_slave_burstcount;    // mm_interconnect_1:address_span_extender_0_windowed_slave_burstcount -> address_span_extender_0:avs_s0_burstcount
	wire  [63:0] mm_interconnect_1_address_span_extender_0_cntl_readdata;                // address_span_extender_0:avs_cntl_readdata -> mm_interconnect_1:address_span_extender_0_cntl_readdata
	wire         mm_interconnect_1_address_span_extender_0_cntl_read;                    // mm_interconnect_1:address_span_extender_0_cntl_read -> address_span_extender_0:avs_cntl_read
	wire   [7:0] mm_interconnect_1_address_span_extender_0_cntl_byteenable;              // mm_interconnect_1:address_span_extender_0_cntl_byteenable -> address_span_extender_0:avs_cntl_byteenable
	wire         mm_interconnect_1_address_span_extender_0_cntl_write;                   // mm_interconnect_1:address_span_extender_0_cntl_write -> address_span_extender_0:avs_cntl_write
	wire  [63:0] mm_interconnect_1_address_span_extender_0_cntl_writedata;               // mm_interconnect_1:address_span_extender_0_cntl_writedata -> address_span_extender_0:avs_cntl_writedata
	wire         mm_interconnect_1_sys_description_rom_s1_chipselect;                    // mm_interconnect_1:sys_description_rom_s1_chipselect -> sys_description_rom:chipselect
	wire  [63:0] mm_interconnect_1_sys_description_rom_s1_readdata;                      // sys_description_rom:readdata -> mm_interconnect_1:sys_description_rom_s1_readdata
	wire         mm_interconnect_1_sys_description_rom_s1_debugaccess;                   // mm_interconnect_1:sys_description_rom_s1_debugaccess -> sys_description_rom:debugaccess
	wire   [8:0] mm_interconnect_1_sys_description_rom_s1_address;                       // mm_interconnect_1:sys_description_rom_s1_address -> sys_description_rom:address
	wire   [7:0] mm_interconnect_1_sys_description_rom_s1_byteenable;                    // mm_interconnect_1:sys_description_rom_s1_byteenable -> sys_description_rom:byteenable
	wire         mm_interconnect_1_sys_description_rom_s1_write;                         // mm_interconnect_1:sys_description_rom_s1_write -> sys_description_rom:write
	wire  [63:0] mm_interconnect_1_sys_description_rom_s1_writedata;                     // mm_interconnect_1:sys_description_rom_s1_writedata -> sys_description_rom:writedata
	wire         mm_interconnect_1_sys_description_rom_s1_clken;                         // mm_interconnect_1:sys_description_rom_s1_clken -> sys_description_rom:clken
	wire  [63:0] mm_interconnect_1_sw_reset_s_readdata;                                  // sw_reset:slave_readdata -> mm_interconnect_1:sw_reset_s_readdata
	wire         mm_interconnect_1_sw_reset_s_waitrequest;                               // sw_reset:slave_waitrequest -> mm_interconnect_1:sw_reset_s_waitrequest
	wire         mm_interconnect_1_sw_reset_s_read;                                      // mm_interconnect_1:sw_reset_s_read -> sw_reset:slave_read
	wire   [7:0] mm_interconnect_1_sw_reset_s_byteenable;                                // mm_interconnect_1:sw_reset_s_byteenable -> sw_reset:slave_byteenable
	wire         mm_interconnect_1_sw_reset_s_write;                                     // mm_interconnect_1:sw_reset_s_write -> sw_reset:slave_write
	wire  [63:0] mm_interconnect_1_sw_reset_s_writedata;                                 // mm_interconnect_1:sw_reset_s_writedata -> sw_reset:slave_writedata
	wire  [31:0] mm_interconnect_1_mem_org_mode_s_readdata;                              // mem_org_mode:slave_readdata -> mm_interconnect_1:mem_org_mode_s_readdata
	wire         mm_interconnect_1_mem_org_mode_s_waitrequest;                           // mem_org_mode:slave_waitrequest -> mm_interconnect_1:mem_org_mode_s_waitrequest
	wire         mm_interconnect_1_mem_org_mode_s_read;                                  // mm_interconnect_1:mem_org_mode_s_read -> mem_org_mode:slave_read
	wire         mm_interconnect_1_mem_org_mode_s_write;                                 // mm_interconnect_1:mem_org_mode_s_write -> mem_org_mode:slave_write
	wire  [31:0] mm_interconnect_1_mem_org_mode_s_writedata;                             // mm_interconnect_1:mem_org_mode_s_writedata -> mem_org_mode:slave_writedata
	wire  [31:0] mm_interconnect_1_version_id_0_s_readdata;                              // version_id_0:slave_readdata -> mm_interconnect_1:version_id_0_s_readdata
	wire         mm_interconnect_1_version_id_0_s_read;                                  // mm_interconnect_1:version_id_0_s_read -> version_id_0:slave_read
	wire  [31:0] mm_interconnect_1_irq_ena_0_s_readdata;                                 // irq_ena_0:slave_readdata -> mm_interconnect_1:irq_ena_0_s_readdata
	wire         mm_interconnect_1_irq_ena_0_s_waitrequest;                              // irq_ena_0:slave_waitrequest -> mm_interconnect_1:irq_ena_0_s_waitrequest
	wire         mm_interconnect_1_irq_ena_0_s_read;                                     // mm_interconnect_1:irq_ena_0_s_read -> irq_ena_0:slave_read
	wire   [3:0] mm_interconnect_1_irq_ena_0_s_byteenable;                               // mm_interconnect_1:irq_ena_0_s_byteenable -> irq_ena_0:slave_byteenable
	wire         mm_interconnect_1_irq_ena_0_s_write;                                    // mm_interconnect_1:irq_ena_0_s_write -> irq_ena_0:slave_write
	wire  [31:0] mm_interconnect_1_irq_ena_0_s_writedata;                                // mm_interconnect_1:irq_ena_0_s_writedata -> irq_ena_0:slave_writedata
	wire         irq_mapper_receiver0_irq;                                               // irq_bridge_0:sender0_irq -> irq_mapper:receiver0_irq
	wire         irq_ena_0_my_irq_in_irq;                                                // irq_mapper:sender_irq -> irq_ena_0:irq
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [irq_ena_0:resetn, kernel_cntrl:reset, mem_org_mode:resetn, mm_interconnect_1:kernel_cntrl_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sys_description_rom:reset, version_id_0:resetn]
	wire         rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [rst_translator:reset_req_in, sys_description_rom:reset_req]
	wire         rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [address_span_extender_0:reset, mm_interconnect_0:address_span_extender_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:address_span_extender_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [mm_interconnect_1:sw_reset_clk_reset_reset_bridge_in_reset_reset, sw_reset:resetn]

	system_acl_iface_acl_kernel_interface_sys_description_rom sys_description_rom (
		.clk         (clk_clk),                                              //   clk1.clk
		.address     (mm_interconnect_1_sys_description_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_sys_description_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_sys_description_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_sys_description_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_sys_description_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_1_sys_description_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_sys_description_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_sys_description_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)                    //       .reset_req
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (30),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) kernel_cra (
		.clk              (kernel_clk_clk),                                //   clk.clk
		.reset            (reset_controller_sw_reset_out_reset),           // reset.reset
		.s0_waitrequest   (mm_interconnect_0_kernel_cra_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_kernel_cra_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_kernel_cra_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_kernel_cra_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_kernel_cra_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_kernel_cra_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_kernel_cra_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_kernel_cra_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_kernel_cra_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_kernel_cra_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (kernel_cra_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (kernel_cra_readdata),                           //      .readdata
		.m0_readdatavalid (kernel_cra_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (kernel_cra_burstcount),                         //      .burstcount
		.m0_writedata     (kernel_cra_writedata),                          //      .writedata
		.m0_address       (kernel_cra_address),                            //      .address
		.m0_write         (kernel_cra_write),                              //      .write
		.m0_read          (kernel_cra_read),                               //      .read
		.m0_byteenable    (kernel_cra_byteenable),                         //      .byteenable
		.m0_debugaccess   (kernel_cra_debugaccess)                         //      .debugaccess
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (30),
		.SLAVE_ADDRESS_WIDTH  (10),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (1),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) address_span_extender_0 (
		.clk                  (kernel_clk_clk),                                                         //           clock.clk
		.reset                (rst_controller_001_reset_out_reset),                                     //           reset.reset
		.avs_s0_address       (mm_interconnect_1_address_span_extender_0_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_1_address_span_extender_0_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_1_address_span_extender_0_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_1_address_span_extender_0_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_1_address_span_extender_0_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_1_address_span_extender_0_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_1_address_span_extender_0_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_1_address_span_extender_0_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_1_address_span_extender_0_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (address_span_extender_0_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (address_span_extender_0_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (address_span_extender_0_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (address_span_extender_0_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (address_span_extender_0_expanded_master_write),                          //                .write
		.avm_m0_writedata     (address_span_extender_0_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (address_span_extender_0_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (address_span_extender_0_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (address_span_extender_0_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_read        (mm_interconnect_1_address_span_extender_0_cntl_read),                    //            cntl.read
		.avs_cntl_readdata    (mm_interconnect_1_address_span_extender_0_cntl_readdata),                //                .readdata
		.avs_cntl_write       (mm_interconnect_1_address_span_extender_0_cntl_write),                   //                .write
		.avs_cntl_writedata   (mm_interconnect_1_address_span_extender_0_cntl_writedata),               //                .writedata
		.avs_cntl_byteenable  (mm_interconnect_1_address_span_extender_0_cntl_byteenable),              //                .byteenable
		.avs_cntl_address     (1'b0)                                                                    //     (terminated)
	);

	sw_reset #(
		.WIDTH             (64),
		.LOG2_RESET_CYCLES (10)
	) sw_reset (
		.clk               (clk_clk),                                  //       clk.clk
		.resetn            (~rst_controller_002_reset_out_reset),      // clk_reset.reset_n
		.slave_write       (mm_interconnect_1_sw_reset_s_write),       //         s.write
		.slave_writedata   (mm_interconnect_1_sw_reset_s_writedata),   //          .writedata
		.slave_byteenable  (mm_interconnect_1_sw_reset_s_byteenable),  //          .byteenable
		.slave_read        (mm_interconnect_1_sw_reset_s_read),        //          .read
		.slave_readdata    (mm_interconnect_1_sw_reset_s_readdata),    //          .readdata
		.slave_waitrequest (mm_interconnect_1_sw_reset_s_waitrequest), //          .waitrequest
		.sw_reset_n_out    (sw_reset_export_reset_n)                   //  sw_reset.reset_n
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (14),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) kernel_cntrl (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (kernel_cntrl_waitrequest),       //    s0.waitrequest
		.s0_readdata      (kernel_cntrl_readdata),          //      .readdata
		.s0_readdatavalid (kernel_cntrl_readdatavalid),     //      .readdatavalid
		.s0_burstcount    (kernel_cntrl_burstcount),        //      .burstcount
		.s0_writedata     (kernel_cntrl_writedata),         //      .writedata
		.s0_address       (kernel_cntrl_address),           //      .address
		.s0_write         (kernel_cntrl_write),             //      .write
		.s0_read          (kernel_cntrl_read),              //      .read
		.s0_byteenable    (kernel_cntrl_byteenable),        //      .byteenable
		.s0_debugaccess   (kernel_cntrl_debugaccess),       //      .debugaccess
		.m0_waitrequest   (kernel_cntrl_m0_waitrequest),    //    m0.waitrequest
		.m0_readdata      (kernel_cntrl_m0_readdata),       //      .readdata
		.m0_readdatavalid (kernel_cntrl_m0_readdatavalid),  //      .readdatavalid
		.m0_burstcount    (kernel_cntrl_m0_burstcount),     //      .burstcount
		.m0_writedata     (kernel_cntrl_m0_writedata),      //      .writedata
		.m0_address       (kernel_cntrl_m0_address),        //      .address
		.m0_write         (kernel_cntrl_m0_write),          //      .write
		.m0_read          (kernel_cntrl_m0_read),           //      .read
		.m0_byteenable    (kernel_cntrl_m0_byteenable),     //      .byteenable
		.m0_debugaccess   (kernel_cntrl_m0_debugaccess)     //      .debugaccess
	);

	mem_org_mode #(
		.WIDTH (32)
	) mem_org_mode (
		.clk                     (clk_clk),                                      //                     clk.clk
		.resetn                  (~rst_controller_reset_out_reset),              //               clk_reset.reset_n
		.slave_write             (mm_interconnect_1_mem_org_mode_s_write),       //                       s.write
		.slave_writedata         (mm_interconnect_1_mem_org_mode_s_writedata),   //                        .writedata
		.slave_read              (mm_interconnect_1_mem_org_mode_s_read),        //                        .read
		.slave_readdata          (mm_interconnect_1_mem_org_mode_s_readdata),    //                        .readdata
		.slave_waitrequest       (mm_interconnect_1_mem_org_mode_s_waitrequest), //                        .waitrequest
		.mem_organization_kernel (acl_bsp_memorg_kernel_mode),                   // mem_organization_kernel.mode
		.mem_organization_host   (acl_bsp_memorg_host_mode)                      //   mem_organization_host.mode
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) irq_bridge_0 (
		.clk          (kernel_clk_clk),                      //          clk.clk
		.receiver_irq (kernel_irq_from_kernel_irq),          // receiver_irq.irq
		.reset        (reset_controller_sw_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_mapper_receiver0_irq),            //  sender0_irq.irq
		.sender1_irq  (),                                    //  (terminated)
		.sender2_irq  (),                                    //  (terminated)
		.sender3_irq  (),                                    //  (terminated)
		.sender4_irq  (),                                    //  (terminated)
		.sender5_irq  (),                                    //  (terminated)
		.sender6_irq  (),                                    //  (terminated)
		.sender7_irq  (),                                    //  (terminated)
		.sender8_irq  (),                                    //  (terminated)
		.sender9_irq  (),                                    //  (terminated)
		.sender10_irq (),                                    //  (terminated)
		.sender11_irq (),                                    //  (terminated)
		.sender12_irq (),                                    //  (terminated)
		.sender13_irq (),                                    //  (terminated)
		.sender14_irq (),                                    //  (terminated)
		.sender15_irq (),                                    //  (terminated)
		.sender16_irq (),                                    //  (terminated)
		.sender17_irq (),                                    //  (terminated)
		.sender18_irq (),                                    //  (terminated)
		.sender19_irq (),                                    //  (terminated)
		.sender20_irq (),                                    //  (terminated)
		.sender21_irq (),                                    //  (terminated)
		.sender22_irq (),                                    //  (terminated)
		.sender23_irq (),                                    //  (terminated)
		.sender24_irq (),                                    //  (terminated)
		.sender25_irq (),                                    //  (terminated)
		.sender26_irq (),                                    //  (terminated)
		.sender27_irq (),                                    //  (terminated)
		.sender28_irq (),                                    //  (terminated)
		.sender29_irq (),                                    //  (terminated)
		.sender30_irq (),                                    //  (terminated)
		.sender31_irq ()                                     //  (terminated)
	);

	version_id #(
		.WIDTH      (32),
		.VERSION_ID (-1598029823)
	) version_id_0 (
		.clk            (clk_clk),                                   //       clk.clk
		.resetn         (~rst_controller_reset_out_reset),           // clk_reset.reset_n
		.slave_read     (mm_interconnect_1_version_id_0_s_read),     //         s.read
		.slave_readdata (mm_interconnect_1_version_id_0_s_readdata)  //          .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_sw (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (~sw_reset_export_reset_n),            // reset_in1.reset
		.clk            (kernel_clk_clk),                      //       clk.clk
		.reset_out      (reset_controller_sw_reset_out_reset), // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	irq_ena irq_ena_0 (
		.clk               (clk_clk),                                   //        clk.clk
		.resetn            (~rst_controller_reset_out_reset),           //  clk_reset.reset_n
		.slave_write       (mm_interconnect_1_irq_ena_0_s_write),       //          s.write
		.slave_writedata   (mm_interconnect_1_irq_ena_0_s_writedata),   //           .writedata
		.slave_byteenable  (mm_interconnect_1_irq_ena_0_s_byteenable),  //           .byteenable
		.slave_read        (mm_interconnect_1_irq_ena_0_s_read),        //           .read
		.slave_readdata    (mm_interconnect_1_irq_ena_0_s_readdata),    //           .readdata
		.slave_waitrequest (mm_interconnect_1_irq_ena_0_s_waitrequest), //           .waitrequest
		.irq               (irq_ena_0_my_irq_in_irq),                   //  my_irq_in.irq
		.irq_out           (kernel_irq_to_host_irq)                     // my_irq_out.irq
	);

	system_acl_iface_acl_kernel_interface_mm_interconnect_0 mm_interconnect_0 (
		.kernel_clk_out_clk_clk                                    (kernel_clk_clk),                                        //                                  kernel_clk_out_clk.clk
		.address_span_extender_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // address_span_extender_0_reset_reset_bridge_in_reset.reset
		.kernel_cra_reset_reset_bridge_in_reset_reset              (reset_controller_sw_reset_out_reset),                   //              kernel_cra_reset_reset_bridge_in_reset.reset
		.address_span_extender_0_expanded_master_address           (address_span_extender_0_expanded_master_address),       //             address_span_extender_0_expanded_master.address
		.address_span_extender_0_expanded_master_waitrequest       (address_span_extender_0_expanded_master_waitrequest),   //                                                    .waitrequest
		.address_span_extender_0_expanded_master_burstcount        (address_span_extender_0_expanded_master_burstcount),    //                                                    .burstcount
		.address_span_extender_0_expanded_master_byteenable        (address_span_extender_0_expanded_master_byteenable),    //                                                    .byteenable
		.address_span_extender_0_expanded_master_read              (address_span_extender_0_expanded_master_read),          //                                                    .read
		.address_span_extender_0_expanded_master_readdata          (address_span_extender_0_expanded_master_readdata),      //                                                    .readdata
		.address_span_extender_0_expanded_master_readdatavalid     (address_span_extender_0_expanded_master_readdatavalid), //                                                    .readdatavalid
		.address_span_extender_0_expanded_master_write             (address_span_extender_0_expanded_master_write),         //                                                    .write
		.address_span_extender_0_expanded_master_writedata         (address_span_extender_0_expanded_master_writedata),     //                                                    .writedata
		.kernel_cra_s0_address                                     (mm_interconnect_0_kernel_cra_s0_address),               //                                       kernel_cra_s0.address
		.kernel_cra_s0_write                                       (mm_interconnect_0_kernel_cra_s0_write),                 //                                                    .write
		.kernel_cra_s0_read                                        (mm_interconnect_0_kernel_cra_s0_read),                  //                                                    .read
		.kernel_cra_s0_readdata                                    (mm_interconnect_0_kernel_cra_s0_readdata),              //                                                    .readdata
		.kernel_cra_s0_writedata                                   (mm_interconnect_0_kernel_cra_s0_writedata),             //                                                    .writedata
		.kernel_cra_s0_burstcount                                  (mm_interconnect_0_kernel_cra_s0_burstcount),            //                                                    .burstcount
		.kernel_cra_s0_byteenable                                  (mm_interconnect_0_kernel_cra_s0_byteenable),            //                                                    .byteenable
		.kernel_cra_s0_readdatavalid                               (mm_interconnect_0_kernel_cra_s0_readdatavalid),         //                                                    .readdatavalid
		.kernel_cra_s0_waitrequest                                 (mm_interconnect_0_kernel_cra_s0_waitrequest),           //                                                    .waitrequest
		.kernel_cra_s0_debugaccess                                 (mm_interconnect_0_kernel_cra_s0_debugaccess)            //                                                    .debugaccess
	);

	system_acl_iface_acl_kernel_interface_mm_interconnect_1 mm_interconnect_1 (
		.clk_reset_clk_clk                                         (clk_clk),                                                                //                                       clk_reset_clk.clk
		.kernel_clk_out_clk_clk                                    (kernel_clk_clk),                                                         //                                  kernel_clk_out_clk.clk
		.address_span_extender_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                     // address_span_extender_0_reset_reset_bridge_in_reset.reset
		.kernel_cntrl_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                         //            kernel_cntrl_reset_reset_bridge_in_reset.reset
		.sw_reset_clk_reset_reset_bridge_in_reset_reset            (rst_controller_002_reset_out_reset),                                     //            sw_reset_clk_reset_reset_bridge_in_reset.reset
		.kernel_cntrl_m0_address                                   (kernel_cntrl_m0_address),                                                //                                     kernel_cntrl_m0.address
		.kernel_cntrl_m0_waitrequest                               (kernel_cntrl_m0_waitrequest),                                            //                                                    .waitrequest
		.kernel_cntrl_m0_burstcount                                (kernel_cntrl_m0_burstcount),                                             //                                                    .burstcount
		.kernel_cntrl_m0_byteenable                                (kernel_cntrl_m0_byteenable),                                             //                                                    .byteenable
		.kernel_cntrl_m0_read                                      (kernel_cntrl_m0_read),                                                   //                                                    .read
		.kernel_cntrl_m0_readdata                                  (kernel_cntrl_m0_readdata),                                               //                                                    .readdata
		.kernel_cntrl_m0_readdatavalid                             (kernel_cntrl_m0_readdatavalid),                                          //                                                    .readdatavalid
		.kernel_cntrl_m0_write                                     (kernel_cntrl_m0_write),                                                  //                                                    .write
		.kernel_cntrl_m0_writedata                                 (kernel_cntrl_m0_writedata),                                              //                                                    .writedata
		.kernel_cntrl_m0_debugaccess                               (kernel_cntrl_m0_debugaccess),                                            //                                                    .debugaccess
		.address_span_extender_0_cntl_write                        (mm_interconnect_1_address_span_extender_0_cntl_write),                   //                        address_span_extender_0_cntl.write
		.address_span_extender_0_cntl_read                         (mm_interconnect_1_address_span_extender_0_cntl_read),                    //                                                    .read
		.address_span_extender_0_cntl_readdata                     (mm_interconnect_1_address_span_extender_0_cntl_readdata),                //                                                    .readdata
		.address_span_extender_0_cntl_writedata                    (mm_interconnect_1_address_span_extender_0_cntl_writedata),               //                                                    .writedata
		.address_span_extender_0_cntl_byteenable                   (mm_interconnect_1_address_span_extender_0_cntl_byteenable),              //                                                    .byteenable
		.address_span_extender_0_windowed_slave_address            (mm_interconnect_1_address_span_extender_0_windowed_slave_address),       //              address_span_extender_0_windowed_slave.address
		.address_span_extender_0_windowed_slave_write              (mm_interconnect_1_address_span_extender_0_windowed_slave_write),         //                                                    .write
		.address_span_extender_0_windowed_slave_read               (mm_interconnect_1_address_span_extender_0_windowed_slave_read),          //                                                    .read
		.address_span_extender_0_windowed_slave_readdata           (mm_interconnect_1_address_span_extender_0_windowed_slave_readdata),      //                                                    .readdata
		.address_span_extender_0_windowed_slave_writedata          (mm_interconnect_1_address_span_extender_0_windowed_slave_writedata),     //                                                    .writedata
		.address_span_extender_0_windowed_slave_burstcount         (mm_interconnect_1_address_span_extender_0_windowed_slave_burstcount),    //                                                    .burstcount
		.address_span_extender_0_windowed_slave_byteenable         (mm_interconnect_1_address_span_extender_0_windowed_slave_byteenable),    //                                                    .byteenable
		.address_span_extender_0_windowed_slave_readdatavalid      (mm_interconnect_1_address_span_extender_0_windowed_slave_readdatavalid), //                                                    .readdatavalid
		.address_span_extender_0_windowed_slave_waitrequest        (mm_interconnect_1_address_span_extender_0_windowed_slave_waitrequest),   //                                                    .waitrequest
		.irq_ena_0_s_write                                         (mm_interconnect_1_irq_ena_0_s_write),                                    //                                         irq_ena_0_s.write
		.irq_ena_0_s_read                                          (mm_interconnect_1_irq_ena_0_s_read),                                     //                                                    .read
		.irq_ena_0_s_readdata                                      (mm_interconnect_1_irq_ena_0_s_readdata),                                 //                                                    .readdata
		.irq_ena_0_s_writedata                                     (mm_interconnect_1_irq_ena_0_s_writedata),                                //                                                    .writedata
		.irq_ena_0_s_byteenable                                    (mm_interconnect_1_irq_ena_0_s_byteenable),                               //                                                    .byteenable
		.irq_ena_0_s_waitrequest                                   (mm_interconnect_1_irq_ena_0_s_waitrequest),                              //                                                    .waitrequest
		.mem_org_mode_s_write                                      (mm_interconnect_1_mem_org_mode_s_write),                                 //                                      mem_org_mode_s.write
		.mem_org_mode_s_read                                       (mm_interconnect_1_mem_org_mode_s_read),                                  //                                                    .read
		.mem_org_mode_s_readdata                                   (mm_interconnect_1_mem_org_mode_s_readdata),                              //                                                    .readdata
		.mem_org_mode_s_writedata                                  (mm_interconnect_1_mem_org_mode_s_writedata),                             //                                                    .writedata
		.mem_org_mode_s_waitrequest                                (mm_interconnect_1_mem_org_mode_s_waitrequest),                           //                                                    .waitrequest
		.sw_reset_s_write                                          (mm_interconnect_1_sw_reset_s_write),                                     //                                          sw_reset_s.write
		.sw_reset_s_read                                           (mm_interconnect_1_sw_reset_s_read),                                      //                                                    .read
		.sw_reset_s_readdata                                       (mm_interconnect_1_sw_reset_s_readdata),                                  //                                                    .readdata
		.sw_reset_s_writedata                                      (mm_interconnect_1_sw_reset_s_writedata),                                 //                                                    .writedata
		.sw_reset_s_byteenable                                     (mm_interconnect_1_sw_reset_s_byteenable),                                //                                                    .byteenable
		.sw_reset_s_waitrequest                                    (mm_interconnect_1_sw_reset_s_waitrequest),                               //                                                    .waitrequest
		.sys_description_rom_s1_address                            (mm_interconnect_1_sys_description_rom_s1_address),                       //                              sys_description_rom_s1.address
		.sys_description_rom_s1_write                              (mm_interconnect_1_sys_description_rom_s1_write),                         //                                                    .write
		.sys_description_rom_s1_readdata                           (mm_interconnect_1_sys_description_rom_s1_readdata),                      //                                                    .readdata
		.sys_description_rom_s1_writedata                          (mm_interconnect_1_sys_description_rom_s1_writedata),                     //                                                    .writedata
		.sys_description_rom_s1_byteenable                         (mm_interconnect_1_sys_description_rom_s1_byteenable),                    //                                                    .byteenable
		.sys_description_rom_s1_chipselect                         (mm_interconnect_1_sys_description_rom_s1_chipselect),                    //                                                    .chipselect
		.sys_description_rom_s1_clken                              (mm_interconnect_1_sys_description_rom_s1_clken),                         //                                                    .clken
		.sys_description_rom_s1_debugaccess                        (mm_interconnect_1_sys_description_rom_s1_debugaccess),                   //                                                    .debugaccess
		.version_id_0_s_read                                       (mm_interconnect_1_version_id_0_s_read),                                  //                                      version_id_0_s.read
		.version_id_0_s_readdata                                   (mm_interconnect_1_version_id_0_s_readdata)                               //                                                    .readdata
	);

	system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (irq_ena_0_my_irq_in_irq)   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (kernel_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (sw_reset_in_reset),                  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign kernel_reset_reset_n = ~reset_controller_sw_reset_out_reset;

endmodule
